module tb;

parameter DWIDTH = 9;
bit		clk=0, rst_n;
logic	enable;

Binary_counter BC(count, clk, rst_n, enable);

always #5 clk = ~clk;

initial 
	begin
	rst_n = 0;
	@(posedge clk); rst_n = 1;
	end
	
initial
	begin
	repeat(20)
		enable = 1;
	$finish;
	end

endmodule