package fifo_package;

typedef enum {STIMULUS, RESET}Pkt_type;
`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "iMonitor.sv"
`include "oMonitor.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"
//`include "top.sv"





endpackage